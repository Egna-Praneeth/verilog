`include "fadder_32.v"

module testbench;
	reg [0:31] in1;
	reg [0:31] in2;
	wire [0:31] sum;
	wire carry;
	
	fadder_32 f1(sum, carry, in1, in2, 1'b0);
	
	initial
		begin
			$monitor(,$time, " in1=%b | in2=%b | sum=%b | carry=%b ", in1, in2, sum, carry);
			#0 in1=32'b00000000000000000000000000000000; in2=32'b00000000000000000000000000000000;
			#3 in1=32'b00000000000000000000000000000001; in2=32'b00000000000000000000000000000000;
			#5 in1=32'b00000000000000000000000000001111; in2=32'b00000000000000000000000000000000;
			#7 in1=32'b00000000000000000000000000000011; in2=32'b00000000000000000000000000000011;
			#9 in1=32'b10000000000000000000000000000000; in2=32'b10000000000000000000000000000000;
			#10 in1=32'b00000000000000000000000000000111; in2=32'b00000000000000000000000000000010;
			#15 $finish;
		end
endmodule